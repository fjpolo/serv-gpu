module barrier_sync #(parameter NUM_CORES = 1) (
    input wire clk,
    input wire rst,
    input wire [NUM_CORES-1:0] core_done, // Signals from cores indicating completion
    output reg all_done                   // Signal indicating all cores are done
);

    reg [NUM_CORES-1:0] done_reg;         // Register to track core completion

    always @(posedge clk or posedge rst) begin
        if (rst) begin
            done_reg <= {NUM_CORES{1'b0}};
            all_done <= 1'b0;
        end else begin
            // Accumulate completion signals
            done_reg <= done_reg | core_done;
            // Check if all cores are done
            if (done_reg == {NUM_CORES{1'b1}})
                all_done <= 1'b1;
        end
    end

endmodule
